// File: tb_ones_count.v

`include "ones_count.v"

module tb_ones_count;

    parameter STEP = 256;

    wire [3:0] count;
    reg [7:0] dat_in;

    ones_count (count, dat_in);

    initial begin
        dat_in = 8'b0;
        for ( k=1; k<STEP; k=k+1 )
            #1 dat_in = dat_in + 1'b1;
    end

    initial begin
        $monitor("At time %4t, dat_in=%b, count=%b",
                    $time, dat_in, count);
    end

endmodule
